library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

--  Uncomment the following lines to use the declarations that are
--  provided for instantiating Xilinx primitive components.
--library UNISIM;
--use UNISIM.VComponents.all;

entity dlx16 is
    Port ( 
    DB: INOUT STD_LOGIC_VECTOR(15 DOWNTO 0);
    AB:BUFFER STD_LOGIC_VECTOR(15 DOWNTO 0);
    MUX: IN STD_LOGIC_VECTOR(0 TO 2);
    CLK,RESET,RUN: IN STD_LOGIC;
    CI:OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
    MWR,MRD,IOW,IOR,MCLK: BUFFER STD_LOGIC;
    PRIX, KRIX: IN STD_LOGIC
    	);
end dlx16;

architecture Behavioral of dlx16 is

	TYPE CMDTYPE IS (T_MOVL, T_MOVH, T_LD, T_ST, T_SLLT, T_MOV, T_SGE, T_ADD, T_SUB, T_AND,
	T_ADDI, T_SUBI, T_ORI, T_BEQZ, T_BNEQ, T_J, T_JAL,T_MOVPC);
	
	FUNCTION DE_INST(INST: STD_LOGIC_VECTOR) RETURN CMDTYPE IS
		BEGIN
		IF(INST = "00000") THEN RETURN T_MOVL;
		ELSIF(INST = "00001") THEN RETURN T_MOVH; 
		ELSIF(INST = "00010") THEN RETURN T_LD;
		ELSIF(INST = "00011") THEN RETURN T_ST;
		ELSIF(INST = "00100") THEN RETURN T_SLLT;
		ELSIF(INST = "00101") THEN RETURN T_MOV;
		ELSIF(INST = "00110") THEN RETURN T_SGE;
		ELSIF(INST = "00111") THEN RETURN T_ADD;
		ELSIF(INST = "01000") THEN RETURN T_SUB;
		ELSIF(INST = "01001") THEN RETURN T_AND;
		ELSIF(INST = "01010") THEN RETURN T_ADDI;
		ELSIF(INST = "01011") THEN RETURN T_SUBI;
		ELSIF(INST = "01100") THEN RETURN T_ORI;
		ELSIF(INST = "01101") THEN RETURN T_BEQZ;
		ELSIF(INST = "01110") THEN RETURN T_BNEQ;
		ELSIF(INST = "01111") THEN RETURN T_J;
		ELSIF(INST = "10000") THEN RETURN T_JAL;
		ELSE RETURN T_MOVPC;
		END IF;
		END FUNCTION;
	
   	SIGNAL R0,R1,R2,R3,R4,R5,R6,R7: STD_LOGIC_VECTOR(15 DOWNTO 0);

-------------------------------

   	FUNCTION GET_REG(REG_NUM: STD_LOGIC_VECTOR) RETURN STD_LOGIC_VECTOR IS
   	BEGIN
   		IF (REG_NUM = "000")THEN 
   			RETURN R0;
   		ELSIF(REG_NUM = "001") THEN
   			RETURN R1;
  	 	ELSIF(REG_NUM = "010") THEN 
   			RETURN R2;
   		ELSIF(REG_NUM = "011") THEN 
   			RETURN R3;
   		ELSIF(REG_NUM = "100") THEN
   			RETURN R4;
   		ELSIF(REG_NUM = "101") THEN
   			RETURN R5;
   		ELSIF(REG_NUM = "110") THEN
   			RETURN R6;
   		ELSE RETURN R7;
   		END IF;
   	END FUNCTION;

  	FUNCTION ISDATA5(INST: CMDTYPE) RETURN BOOLEAN IS
   	BEGIN
   			IF (INST = T_LD OR INST = T_ST OR INST = T_MOV) THEN
   				RETURN TRUE;
   			ELSE RETURN FALSE;
   			END IF;
   	END FUNCTION;

   	FUNCTION ISDATA8(INST: CMDTYPE) RETURN BOOLEAN IS
   	BEGIN
   			IF (INST = T_ADDI OR INST = T_SUBI OR INST = T_ORI OR INST = T_BEQZ OR INST = T_BNEQ OR INST = T_MOVPC) THEN
   				RETURN TRUE;
   			ELSE RETURN FALSE;
   			END IF;
   	END FUNCTION;

   	FUNCTION ISJMP(INST: CMDTYPE) RETURN BOOLEAN IS
   	BEGIN
   			IF (INST = T_J OR INST = T_JAL) THEN
   				RETURN TRUE;
   			ELSE RETURN FALSE;
   			END IF;
   	END FUNCTION;

   	FUNCTION USEA(INST: CMDTYPE) RETURN BOOLEAN IS
   	BEGIN
   			IF(INST = T_LD OR INST = T_ST OR INST = T_SLLI OR INST = T_MOV OR INST = T_SGE  OR INST = T_ADD OR INST = T_SUB OR INST = T_AND 
        	OR INST = T_ADDI OR INST = T_SUBI OR INST = T_ORI OR INST = T_BEQZ OR INST = T_BNEQ OR INST = T_MOVPC OR INST = T_MOVL OR INST = T_MOVH)
   				THEN RETURN TRUE;
   			ELSE RETURN FALSE;
   			END IF;
   	END FUNCTION;

   	FUNCTION USEB(INST: CMDTYPE) RETURN BOOLEAN IS
   	BEGIN 
   			IF(INST = T_SGE OR INST = T_ADD OR INST = T_SUB OR INST = T_AND)
   				THEN RETURN TRUE;
   			ELSE RETURN FALSE;
   			END IF;
   	END FUNCTION;

   	FUNCTION USEW(INST: CMDTYPE) RETURN BOOLEAN IS
   	BEGIN
   			IF(INST = T_MOVL OR INST = T_MOVH OR INST = T_LD OR INST = T_SLLT OR INST = T_MOV 
   				OR INST = T_SGE OR INST = T_ADD OR INST = T_SUB OR INST = T_ADDI OR INST = SUNBI
   				OR INST = ORI OR INST = T_JAL)
   				THEN RETURN TRUE;
   			ELSE RETURN FALSE;
   			END IF;
   	END FUNCTION;

   	FUNCTION EXTO16(NUM:STD_LOGIC_VECTOR; LEN: INTEGER) RETURN STD_LOGIC_VECTOR IS
   		VARIABLE RES : STD_LOGIC_VECTOR(15 DOWNTO 0);
   		VARIABLE I : INTEGER;
   	BEGIN
   		FOR I IN LEN TO 15 LOOP
   			RES(I) := NUM(LEN-1);
   		END LOOP;
   		RES(LEN-1 DOWNTO 0) := NUM;
   		RETURN RES;
   	END FUNCTION;

   	FUNCTION REG_W1(INST: CMDTYPE) RETURN BOOLEAN IS
   	BEGIN 
   		IF (INST = T_MOVL OR INST = T_MOVH OR INST = T_ADDI OR INST = T_SUBI OR INST = T_ORI)
   			THEN RETURN TRUE;
   		ELSE RETURN FALSE;
   		END IF;
   	END FUNCTION;

   	FUNCTION REG_W2(INST: CMDTYPE) RETURN BOOLEAN IS
   	BEGIN 
   		IF (INST = T_MOV OR INST = T_SLLT OR INST = T_LD)
   			THEN RETURN TRUE;
   		ELSE RETURN FALSE;
   		END IF;
   	END FUNCTION;

   	FUNCTION REG_W3(INST: CMDTYPE) RETURN BOOLEAN IS
   	BEGIN 
   		IF (INST = T_SGE OR INST = T_AND OR INST = T_SUB OR INST = T_ADD)
   			THEN RETURN TRUE;
   		ELSE RETURN FALSE;
   		END IF;
   	END FUNCTION;

   	SIGNAL ID_INS, EX_INS,ME_INS, WB_INS: CMDTYPE;
   	SIGNAL ID_REGA, ID_REGB, EX_REGA, EX_REGB, EX_REGW, ME_REGB, ME_REGW,WB_REGW: STD_LOGIC_VECTOR(2 DOWNTO 0);
   	SIGNAL ID_USEA, ID_USEB, EX_USEA, EX_USEB, EX_USEW, ME_USEW, WB_USEW: STD_LOGIC;
   	SIGNAL ME_W_DATA, WB_W_DATA: STD_LOGIC_VECTOR(15 DOWNTO 0);
   	SIGNAL PC: STD_LOGIC_VECTOR(15 DOWNTO 0);
   	SIGNAL MUXAB: STD_LOGIC_VECTOR(15 DOWNTO 0);
   	SIGNAL STALL, BUBBLE: STD_LOGIC_VECTOR(0 TO 4);
   	SIGNAL OB, WRE: STD_LOGIC;
   	SIGNAL IR_ID, IR_EX, IR_ME, IR_WB: STD_LOGIC_VECTOR(15 DOWNTO 0);
   	SIGNAL PC_ID, PC_EX, PC_ME, PC_WB: STD_LOGIC_VECTOR(15 DOWNTO 0);
   	SIGNAL ID_IMM, EX_A, EX_B, EX_IMM: STD_LOGIC_VECTOR(15 DOWNTO 0);
   	
   	SIGNAL BUF_STALL, BUF_BUBBLE: STD_LOGIC_VECTOR(0 TO 4);
   	SIGNAL BUF_PC: STD_LOGIC_VECTOR(15 DOWNTO 0);
   	SIGNAL BUF_ID_REGA, BUF_ID_REGB: STD_LOGIC_VECTOR(15 DOWNTO 0);
   	SIGNAL BUF_ID_DATAA, BUF_ID_DATAB: STD_LOGIC_VECTOR(15 DOWNTO 0);
   	SIGNAL BUF_ID_OUT: STD_LOGIC_VECTOR(15 DOWNTO 0);
   	SIGNAL BUF_ID_MIS: STD_LOGIC;
   	SIGNAL BUF_EX_DATAA, BUF_EX_DATAB: STD_LOGIC_VECTOR(15 DOWNTO 0);
   	SIGNAL BUF_EX_MUXA, BUF_EX_MUXB: STD_LOGIC_VECTOR(15 DOWNTO 0);
   	SIGNAL BUF_EX_OUT: STD_LOGIC_VECTOR(15 DOWNTO 0);
   	SIGNAL BUF_EX_TMP: STD_LOGIC_VECTOR(15 DOWNTO 0);
   	SIGNAL BUF_ME_DATA: STD_LOGIC_VECTOR(15 DOWNTO 0);
   	SIGNAL BUF_ME_B: STD_LOGIC_VECTOR(15 DOWNTO 0);
   	SIGNAL ME_B, ME_OUT: STD_LOGIC_VECTOR(15 DOWNTO 0);
   	SIGNAL WB_MEM_DATA,WB_OUT: STD_LOGIC_VECTOR(15 DOWNTO 0);

   	SIGNAL MIS: BOOLEAN;
   	SIGNAL LOADUSEH: BOOLEAN;
   	SIGNAL STR: BOOLEAN;


BEGIN
	
	PROCESS(MCLK,CLK) BEGIN
		IF RUN = '0' OR RESET = '0' THEN MCLK <= '0';
		ELSIF CLK'EVENT AND CLK = '0' THEN MCLK <= NOT MCLK;
		END IF;
	END PROCESS;

	ID_INS <= DE_INST(IR_ID(15 DOWNTO 11));
	EX_INS <= DE_INST(EX_ID(15 DOWNTO 11));
	ME_INS <= DE_INST(ME_ID(15 DOWNTO 11));
	WB_INS <= DE_INST(WB_ID(15 DOWNTO 11));

---ID

	ID_REGA <= IR_ID(10 DOWNTO 8);
	ID_REGB <= IR_ID(7 DOWNTO 5);
	ID_USEA <= '1' WHEN USEA(ID_INS) ELSE '0';
	ID_USEB <= '1' WHEN USEB(ID_INS) ELSE '0'; 

	ID_IMM <= EXTO16(IR_ID(10 DOWNTO 0),11) WHEN ISJMP(ID_INS) ELSE
				EXTO16(IR_ID(7 DOWNTO 0), 8) WHEN ISDATA8(ID_INS) ELSE
				EXTO16(IR_ID(4 DOWNTO 0), 5) WHEN ISDATA5(ID_INS) ELSE
				"00000000" & IR_ID(7 DOWNTO 0) WHEN ID_INS = T_MOVL ELSE
				IR_ID(7 DOWNTO 0) & "00000000" WHEN ID_INS = T_MOVH ELSE
				"00000000000" & IR_ID(4 DOWNTO 0);

---EX

	EX_REGA <= IR_EX(10 DOWNTO 8);
	EX_REGB <= IR_EX(7 DOWNTO 5);
	EX_USEA <= '1' WHEN USEA(EX_INS) ELSE '0';
	EX_USEB <= '1' WHEN USEB(EX_INS) ELSE '0';
	EX_USEW <= '1' WHEN USEW(EX_INS) ELSE '0';

	EX_IMM <= EXTO16(IR_EX(10 DOWNTO 0),11) WHEN ISJMP(EX_INS) ELSE
				EXTO16(IR_EX(7 DOWNTO 0),8) WHEN ISDATA8(EX_INS) ELSE
				EXTO16(IR_EX(4 DOWNTO 0),5) WHEN ISDATA5(EX_INS) ELSE
				"00000000" & IR_EX(7 DOWNTO 0) WHEN EX_INS = T_MOVL ELSE
				IR_EX(7 DOWNTO 0) & "00000000" WHEN EX_INS = T_MOVH ELSE
				"00000000000" & IR_EX(4 DOWNTO 0);

	EX_REGW <= IR_EX(10 DOWNTO 8) WHEN REG_W1(EX_INS) ELSE
			IR_EX(7 DOWNTO 5) WHEN REG_W2(EX_INS) ELSE
			IR_EX(4 DOWNTO 2) WHEN REG_W3(EX_INS) ELSE
			"111";

---MEM

	ME_REGB <= IR_ME(7 DOWNTO 5);
	ME_USEW <= '1' WHEN USEW(ME_INS) ELSE '0';

	ME_REGW <= IR_ME(10 DOWNTO 8) WHEN REG_W1(ME_INS) ELSE
			IR_ME(7 DOWNTO 5) WHEN REG_W2(ME_INS) ELSE
			IR_ME(4 DOWNTO 2) WHEN REG_W3(ME_INS) ELSE
			"111";

	ME_W_DATA <= BUF_ME_DATA WHEN ME_INS = T_LD ELSE
				PC_ME WHEN ME_INS = T_JAL ELSE ME_OUT;

---WB
	
	WB_USEW <= '1' WHEN USEW(WB_INS) ELSE '0';

	WB_REGW <= IR_RB(10 DOWNTO 8) WHEN IR_WB(15 DOWNTO 11) = "00000" OR
				IR_WB(15 DOWNTO 11) = "00001" OR IR_WB(15 DOWNTO 11) = "01010" OR
				IR_WB(15 DOWNTO 11) = "01011" OR IR_WB(15 DOWNTO 11) = "01100" ELSE
				IR_WB(7 DOWNTO 5) WHEN REG_W2(WB_INS) ELSE
				IR_WB(4 DOWNTO 2) WHEN REG_W3(WB_INS) ELSE
				"111";

	WB_W_DATA <= WB_MEM_DATA WHEN WB_INS = T_LD ELSE
				PC_WB WHEN WB_INS = T_JAL ELSE
				WB_OUT;

---AB

	MUXAB <= PC WHEN BUBBLE(0) = '1' ELSE ME_OUT;
	AB <= MUXAB;

	BUF_ME_DATA <= DB WHEN (AB(15) = '0' OR AB = "1000000000000001") AND ME_INS = T_LD AND BUBBLE(3) = '1' ELSE
				"000000000000000" & KRIX WHEN AB(15) = '1' AND AB(2) = '1' ELSE
				"000000000000000" & PRIX;

---DB

	OB <= '0' WHEN BUBBLE(3) = '1' AND ME_INS = T_ST ELSE '1';
	DB <= BUF_ME_B WHEN OB = '0' ELSE "ZZZZZZZZZZZZZZZZ";

---RD/WB

	MRD <= '0' WHEN BUBBLE(0) = '1' OR (bubble(3) = '1' AND ME_INS = T_LD and AB(15) = '0') ELSE '1';
    MWR <= '0' WHEN BUBBLE(3) = '1' AND ME_INS = T_ST AND AB(15) = '0' AND MCLK = '1' ELSE '1';

    IOR <= '0' WHEN bubble(3) = '1' AND ME_CMD = T_LD AND AB(15) = '1' AND AB(0) = '1' ELSE '1';
    IOW <= '0' WHEN bubble(3) = '1' AND ME_CMD = T_ST and AB(15) = '1' and AB(1) = '1' and MCLK = '1' else '1';

	WRE <= '1' WHEN bubble(4) = '0' OR WB_CMD = T_ST OR WB_CMD = T_BEQZ OR WB_CMD = T_BNEQ 
			OR WB_CMD = T_J OR WB_CMD = T_MOVPC ELSE '0';


	MIS <= TRUE WHEN BUBBLE(1) = '1' AND BUF_ID_MIS = '1' ELSE FALSE;
	LOADUSEH <= TRUE WHEN BUBBLE(2) = '1' AND BUBBLE(1) = '1' AND EX_INS = T_LD
					AND ((ID_USEA = '1' AND ID_REGA = EX_REGW) OR (ID_USEB = '1' AND ID_REGB = EX_REGW)) ELSE FALSE;
	STR <= TRUE WHEN BUBBLE(2) = '1' AND (EX_INS = T_LD OR EX_INS = T_ST) ELSE FALSE;

	BUF_STALL <= "00111" WHEN LOADUSEH ELSE "11111";
	BUF_BUBBLE <= "000" & BUBBLE(2) & BUBBLE(3) WHEN MIS AND LOADUSEH AND STR ELSE
				'0' & BUBBLE(0) & '0' & BUBBLE(2) & BUBBLE(3) WHEN LOADUSEH AND STR ELSE
				'1' & BUBBLE(0) & '0' & BUBBLE(2) & BUBBLE(3) WHEN LOADUSEH ELSE
				'0' & BUBBLE(0) & BUBBLE(1) & BUBBLE(2) & BUBBLE(3) WHEN STR ELSE
				"10" & BUBBLE(1) & BUBBLE(2) & BUBBLE(3) WHEN MIS ELSE
				"100" & BUBBLE(2) & BUBBLE(3) & WHEN LOADUSEH AND MIS ELSE
				"00" & BUBBLE(1) & BUBBLE(2) & BUBBLE(3) WHEN STR AND MIS ELSE
				'1' & BUBBLE(0) & BUBBLE(1) & BUBBLE(2) & BUBBLE(3);

----------------

	BUF_PC <= BUF_ID_OUT WHEN BUBBLE(1) = '1' AND BUF_ID_MIS = '1' ELSE
			PC + 1 WHEN BUBBLE(0) = '1' ELSE PC;

----------------

	BUF_ID_REGA <= DE_INST(ID_REGA);
	BUF_ID_REGB <= DE_INST(ID_REGB);

	BUF_ID_DATAA <= WB_W_DATA WHEN BUBBLE(4) = '1' AND WB_USEW = '1' AND WB_REGW = ID_REGA ELSE
					ME_W_DATA WHEN BUBBLE(3) = '1' AND ME_USEW = '1' AND ME_REGW = ID_REGA ELSE
					BUF_EX_OUT WHEN BUBBLW(2) = '1' AND EX_USEW = '1' AND EX_REGW = ID_REGA ELSE
					BUF_ID_REGA;

	BUF_ID_DATAB <= WB_W_DATA WHEN BUBBLE(4) = '1' AND WB_USEW = '1' AND WB_REGW = ID_REGB ELSE
					ME_W_DATA WHEN BUBBLE(3) = '1' AND ME_USEW = '1' AND ME_REGW = ID_REGB ELSE
					BUF_EX_OUT WHEN BUBBLW(2) = '1' AND EX_USEW = '1' AND EX_REGW = ID_REGB ELSE
					BUF_ID_REGB;

	BUF_ID_MIS <= '1' WHEN ID_INS = T_J OR ID_INS = T_JAL OR ID_INS = T_MOVPC ELSE
					'1' WHEN BUF_BUBBLE(2) = '1' AND ((ID_INS = T_BEQZ AND BUF_ID_DATAA = "0000000000000000") OR (ID_INS = T_BNEQ AND BUF_ID_DATAA /= "0000000000000000")) ELSE
					'0';

	BUF_ID_OUT <= ID_PC + ID_IMM WHEN ID_INS /= T_MOVPC ELSE BUF_ID_DATAA;

----------------

	BUF_EX_DATAA <= WB_W_DATA WHEN BUBBLE(4) = '1' AND WB_USEW = '1' AND WB_REGW = EX_REGA ELSE
					ME_W_DATA WHEN BUBBLE(3) = '1' AND ME_USEW = '1' AND ME_REGW = EX_REGA ELSE
					EX_A;

	BUF_EX_DATAB <= WB_W_DATA WHEN BUBBLE(4) = '1' AND WB_USEW = '1' AND WB_REGW = EX_REGB ELSE
					ME_W_DATA WHEN BUBBLE(3) = '1' AND ME_USEW = '1' AND ME_REGW = EX_REGB ELSE
					EX_B;

	BUF_EX_MUXA <= BUF_EX_DATAA(15 DOWNTO 8) & "00000000" WHEN EX_INS = T_MOVL ELSE
					"00000000" & BUF_EX_DATAA(7 DOWNTO 0) WHEN EX_INS = T_MOVH ELSE
					BUF_EX_DATAA;

	BUF_EX_MUXB <= BUF_EX_DATAB WHEN EX_INS = T_SGE OR EX_INS = T_ADD OR EX_INS = T_SUB OR EX_INS = T_AND ELSE
					EX_IMM;

-------ALU------

	BUF_EX_TMP <= BUF_EX_MUXA - BUF_EX_MUXB;

	BUF_EX_OUT <= BUF_EX_MUXA - BUF_EX_MUXB WHEN EX_INS = T_SUB OR EX_INS = T_SUBI ELSE
					BUF_EX_MUXA AND BUF_EX_MUXB WHEN EX_INS = T_AND ELSE
					BUF_EX_MUXA OR BUF_EX_MUXB WHEN EX_INS = T_ORI ELSE
					TO_STDLOGICVECTOR(TO_BITVECTOR(BUF_EX_MUXA) SLL CONV_INTEGER(BUF_EX_MUXB)) WHEN EX_INS = T_SLLI ELSE
					"0000000000000001" WHEN BUF_EX_TMP(15) = '0' AND EX_INS = T_SGE ELSE
					"0000000000000000" WHEN BUF_EX_TMP(15) = '1' AND EX_INS = T_SGE ELSE
					BUF_EX_MUXA + BUF_EX_MUXB;

----------------

	BUF_ME_B <= WB_W_DATA WHEN BUBBLE(4) = '1' AND WB_USEW = '1' AND WB_REGW = ME_REGB ELSE
				ME_B;

----------------

	PROCESS(MCLK) BEGIN
		IF MCLK'EVENT AND MCLK = '1' THEN 
			IF BUBBLE(4) = '1' AND WRE = '0' THEN 
				IF WB_REGW = "000" THEN R0 <= WB_W_DATA;
				ELSIF WB_REGW = "001" THEN R1 <= WB_W_DATA;
				ELSIF WB_REGW = "010" THEN R2 <= WB_W_DATA;
				ELSIF WB_REGW = "011" THEN R3 <= WB_W_DATA;
				ELSIF WB_REGW = "100" THEN R4 <= WB_W_DATA;
				ELSIF WB_REGW = "101" THEN R5 <= WB_W_DATA;
				ELSIF WB_REGW = "110" THEN R6 <= WB_W_DATA;
				ELSE R7 <= WB_W_DATA;
				END IF;
			END IF;
		END IF;
	END PROCESS;

	PROCESS(MCLK, RUN, RESET) BEGIN
		IF RUN = '0' OR RESET = '0' THEN 
			PC <= "0000000000000000";
			BUBBLE <= "10000";
			STALL <= "11111";
			IR_ID <= "1111111111111111";
			IR_EX <= "1111111111111111";
			IR_ME <= "1111111111111111";
			IR_WB <= "1111111111111111";

		ELSIF MCLK'EVENT AND MCLK = '0' THEN
			IF BUF_STALL(4) = '1' THEN
				IR_WB <= IR_ME;
				PC_WB <= PC_ME;
				WB_OUT <= ME_OUT;
				WB_MEM_DATA <= BUF_ME_DATA;
			END IF;

			IF BUF_STALL(3) = '1' THEN
				IR_ME <= IR_EX;
				PC_ME <= PC_EX;
				ME_OUT <= BUF_EX_OUT;
				ME_B <= BUF_EX_DATAB;
			END IF;

			IF BUF_STALL(2) = '1' THEN
				IR_EX <= IR_ID;
				PC_EX <= PC_ID;
				EX_A <= BUF_ID_DATAA;
				EX_B <= BUF_ID_DATAB;
			END IF;

			IF BUF_STALL(1) = '1' THEN
				PC_ID <= PC + 1;
				IR_ID <= DB;
			END IF;

			IF BUF_STALL(0) = '1' THEN
				PC <= BUF_PC;
			END IF;

			STALL <= BUF_STALL;
			BUBBLE <= BUF_BUBBLE;

		END IF;

	END PROCESS;

	CI(31 DOWNTO 16) <= IR_ID WHEN MUX = "000" ELSE
						IR_EX WHEN MUX = "001" ELSE
						IR_ME WHEN MUX = "010" ELSE
						IR_WB WHEN MUX = "011" ELSE
						R4 WHEN MUX = "100" ELSE
						R5 WHEN MUX = "101" ELSE
						R6 WHEN MUX = "110" ELSE
						R7;

	CI(15 DOWNTO 0) <=  PC WHEN MUX = "000" ELSE
						ME_B WHEN MUX = "001" ELSE
						STALL & BUBBLE & WRE & PRIX & KRIX & BUF_ID_MIS & OB & '0' WHEN MUX = "010" ELSE
						WB_MEM_DATA WHEN MUX = "011" ELSE
						R0 WHEN MUX = "100" ELSE
						R1 WHEN MUX = "101" ELSE
						R2 WHEN MUX = "110" ELSE
						R3;

end Behavioral;
